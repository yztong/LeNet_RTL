//==================================================================================================
//  Filename      : w5_rom.v
//  Created On    : 2018-01-07 22:27:49
//  Last Modified : 2018-03-21 15:10:42
//  Revision      : 
//  Author        : YzTong
//  Company       : UESTC
//  Email         : yztong1994@gmail.com
//
//  Description   : 
//
//
//==================================================================================================
module w5_rom(/*autoport*/
//output
      w5_1_rdata,
      w5_2_rdata,
      w5_3_rdata,
      w5_4_rdata,
      w5_5_rdata,
      w5_6_rdata,
      w5_7_rdata,
      w5_8_rdata,
      w5_9_rdata,
      w5_10_rdata,
      w5_11_rdata,
      w5_12_rdata,
      w5_13_rdata,
      w5_14_rdata,
      w5_15_rdata,
      w5_16_rdata,
      w5_17_rdata,
      w5_18_rdata,
      w5_19_rdata,
      w5_20_rdata,
      w5_21_rdata,
      w5_22_rdata,
      w5_23_rdata,
      w5_24_rdata,
      w5_25_rdata,
      w5_26_rdata,
      w5_27_rdata,
      w5_28_rdata,
      w5_29_rdata,
      w5_30_rdata,
      w5_31_rdata,
      w5_32_rdata,
      w5_33_rdata,
      w5_34_rdata,
      w5_35_rdata,
      w5_36_rdata,
      w5_37_rdata,
      w5_38_rdata,
      w5_39_rdata,
      w5_40_rdata,
      w5_41_rdata,
      w5_42_rdata,
      w5_43_rdata,
      w5_44_rdata,
      w5_45_rdata,
      w5_46_rdata,
      w5_47_rdata,
      w5_48_rdata,
      w5_49_rdata,
      w5_50_rdata,
      w5_51_rdata,
      w5_52_rdata,
      w5_53_rdata,
      w5_54_rdata,
      w5_55_rdata,
      w5_56_rdata,
      w5_57_rdata,
      w5_58_rdata,
      w5_59_rdata,
      w5_60_rdata,
      w5_61_rdata,
      w5_62_rdata,
      w5_63_rdata,
      w5_64_rdata,
      w5_65_rdata,
      w5_66_rdata,
      w5_67_rdata,
      w5_68_rdata,
      w5_69_rdata,
      w5_70_rdata,
      w5_71_rdata,
      w5_72_rdata,
      w5_73_rdata,
      w5_74_rdata,
      w5_75_rdata,
      w5_76_rdata,
      w5_77_rdata,
      w5_78_rdata,
      w5_79_rdata,
      w5_80_rdata,
      w5_81_rdata,
      w5_82_rdata,
      w5_83_rdata,
      w5_84_rdata,
      w5_85_rdata,
      w5_86_rdata,
      w5_87_rdata,
      w5_88_rdata,
      w5_89_rdata,
      w5_90_rdata,
      w5_91_rdata,
      w5_92_rdata,
      w5_93_rdata,
      w5_94_rdata,
      w5_95_rdata,
      w5_96_rdata,
      w5_97_rdata,
      w5_98_rdata,
      w5_99_rdata,
      w5_100_rdata,
      w5_101_rdata,
      w5_102_rdata,
      w5_103_rdata,
      w5_104_rdata,
      w5_105_rdata,
      w5_106_rdata,
      w5_107_rdata,
      w5_108_rdata,
      w5_109_rdata,
      w5_110_rdata,
      w5_111_rdata,
      w5_112_rdata,
      w5_113_rdata,
      w5_114_rdata,
      w5_115_rdata,
      w5_116_rdata,
      w5_117_rdata,
      w5_118_rdata,
      w5_119_rdata,
      w5_120_rdata,
//input
      clk,
      w5_raddr);
	
	input clk;
	input [8:0] w5_raddr;
	output[7:0] w5_1_rdata;	
	output[7:0] w5_2_rdata;
	output[7:0] w5_3_rdata;
	output[7:0] w5_4_rdata;
	output[7:0] w5_5_rdata;
	output[7:0] w5_6_rdata;
	output[7:0] w5_7_rdata;
	output[7:0] w5_8_rdata;
	output[7:0] w5_9_rdata;
	output[7:0] w5_10_rdata;
	output[7:0] w5_11_rdata;
	output[7:0] w5_12_rdata;
	output[7:0] w5_13_rdata;
	output[7:0] w5_14_rdata;
	output[7:0] w5_15_rdata;
	output[7:0] w5_16_rdata;
	output[7:0] w5_17_rdata;
	output[7:0] w5_18_rdata;
	output[7:0] w5_19_rdata;
	output[7:0] w5_20_rdata;
	output[7:0] w5_21_rdata;
	output[7:0] w5_22_rdata;
	output[7:0] w5_23_rdata;
	output[7:0] w5_24_rdata;
	output[7:0] w5_25_rdata;
	output[7:0] w5_26_rdata;
	output[7:0] w5_27_rdata;
	output[7:0] w5_28_rdata;
	output[7:0] w5_29_rdata;
	output[7:0] w5_30_rdata;
	output[7:0] w5_31_rdata;
	output[7:0] w5_32_rdata;
	output[7:0] w5_33_rdata;
	output[7:0] w5_34_rdata;
	output[7:0] w5_35_rdata;
	output[7:0] w5_36_rdata;
	output[7:0] w5_37_rdata;
	output[7:0] w5_38_rdata;
	output[7:0] w5_39_rdata;
	output[7:0] w5_40_rdata;
	output[7:0] w5_41_rdata;
	output[7:0] w5_42_rdata;
	output[7:0] w5_43_rdata;
	output[7:0] w5_44_rdata;
	output[7:0] w5_45_rdata;
	output[7:0] w5_46_rdata;
	output[7:0] w5_47_rdata;
	output[7:0] w5_48_rdata;
	output[7:0] w5_49_rdata;
	output[7:0] w5_50_rdata;
	output[7:0] w5_51_rdata;
	output[7:0] w5_52_rdata;
	output[7:0] w5_53_rdata;
	output[7:0] w5_54_rdata;
	output[7:0] w5_55_rdata;
	output[7:0] w5_56_rdata;
	output[7:0] w5_57_rdata;
	output[7:0] w5_58_rdata;
	output[7:0] w5_59_rdata;
	output[7:0] w5_60_rdata;
	output[7:0] w5_61_rdata;
	output[7:0] w5_62_rdata;
	output[7:0] w5_63_rdata;
	output[7:0] w5_64_rdata;
	output[7:0] w5_65_rdata;
	output[7:0] w5_66_rdata;
	output[7:0] w5_67_rdata;
	output[7:0] w5_68_rdata;
	output[7:0] w5_69_rdata;
	output[7:0] w5_70_rdata;
	output[7:0] w5_71_rdata;
	output[7:0] w5_72_rdata;
	output[7:0] w5_73_rdata;
	output[7:0] w5_74_rdata;
	output[7:0] w5_75_rdata;
	output[7:0] w5_76_rdata;
	output[7:0] w5_77_rdata;
	output[7:0] w5_78_rdata;
	output[7:0] w5_79_rdata;
	output[7:0] w5_80_rdata;
	output[7:0] w5_81_rdata;
	output[7:0] w5_82_rdata;
	output[7:0] w5_83_rdata;
	output[7:0] w5_84_rdata;
	output[7:0] w5_85_rdata;
	output[7:0] w5_86_rdata;
	output[7:0] w5_87_rdata;
	output[7:0] w5_88_rdata;
	output[7:0] w5_89_rdata;
	output[7:0] w5_90_rdata;
	output[7:0] w5_91_rdata;
	output[7:0] w5_92_rdata;
	output[7:0] w5_93_rdata;
	output[7:0] w5_94_rdata;
	output[7:0] w5_95_rdata;
	output[7:0] w5_96_rdata;
	output[7:0] w5_97_rdata;
	output[7:0] w5_98_rdata;
	output[7:0] w5_99_rdata;
	output[7:0] w5_100_rdata;
	output[7:0] w5_101_rdata;
	output[7:0] w5_102_rdata;
	output[7:0] w5_103_rdata;
	output[7:0] w5_104_rdata;
	output[7:0] w5_105_rdata;
	output[7:0] w5_106_rdata;
	output[7:0] w5_107_rdata;
	output[7:0] w5_108_rdata;
	output[7:0] w5_109_rdata;
	output[7:0] w5_110_rdata;
	output[7:0] w5_111_rdata;
	output[7:0] w5_112_rdata;
	output[7:0] w5_113_rdata;
	output[7:0] w5_114_rdata;
	output[7:0] w5_115_rdata;
	output[7:0] w5_116_rdata;
	output[7:0] w5_117_rdata;
	output[7:0] w5_118_rdata;
	output[7:0] w5_119_rdata;
	output[7:0] w5_120_rdata;


  wire [959:0] w5_rdata;
  blk_mem_gen_w5_rom w5_rom (
    .clka(clk),    // input clka
    .addra(w5_raddr),  // input [8 : 0] addra
    .douta(w5_rdata)  // output [959 : 0] douta
  );

  assign w5_1_rdata = w5_rdata[7:0];
  assign w5_2_rdata = w5_rdata[15:8];
  assign w5_3_rdata = w5_rdata[23:16];
  assign w5_4_rdata = w5_rdata[31:24];
  assign w5_5_rdata = w5_rdata[39:32];
  assign w5_6_rdata = w5_rdata[47:40];
  assign w5_7_rdata = w5_rdata[55:48];
  assign w5_8_rdata = w5_rdata[63:56];
  assign w5_9_rdata = w5_rdata[71:64];
  assign w5_10_rdata = w5_rdata[79:72];
  assign w5_11_rdata = w5_rdata[87:80];
  assign w5_12_rdata = w5_rdata[95:88];
  assign w5_13_rdata = w5_rdata[103:96];
  assign w5_14_rdata = w5_rdata[111:104];
  assign w5_15_rdata = w5_rdata[119:112];
  assign w5_16_rdata = w5_rdata[127:120];
  assign w5_17_rdata = w5_rdata[135:128];
  assign w5_18_rdata = w5_rdata[143:136];
  assign w5_19_rdata = w5_rdata[151:144];
  assign w5_20_rdata = w5_rdata[159:152];
  assign w5_21_rdata = w5_rdata[167:160];
  assign w5_22_rdata = w5_rdata[175:168];
  assign w5_23_rdata = w5_rdata[183:176];
  assign w5_24_rdata = w5_rdata[191:184];
  assign w5_25_rdata = w5_rdata[199:192];
  assign w5_26_rdata = w5_rdata[207:200];
  assign w5_27_rdata = w5_rdata[215:208];
  assign w5_28_rdata = w5_rdata[223:216];
  assign w5_29_rdata = w5_rdata[231:224];
  assign w5_30_rdata = w5_rdata[239:232];
  assign w5_31_rdata = w5_rdata[247:240];
  assign w5_32_rdata = w5_rdata[255:248];
  assign w5_33_rdata = w5_rdata[263:256];
  assign w5_34_rdata = w5_rdata[271:264];
  assign w5_35_rdata = w5_rdata[279:272];
  assign w5_36_rdata = w5_rdata[287:280];
  assign w5_37_rdata = w5_rdata[295:288];
  assign w5_38_rdata = w5_rdata[303:296];
  assign w5_39_rdata = w5_rdata[311:304];
  assign w5_40_rdata = w5_rdata[319:312];
  assign w5_41_rdata = w5_rdata[327:320];
  assign w5_42_rdata = w5_rdata[335:328];
  assign w5_43_rdata = w5_rdata[343:336];
  assign w5_44_rdata = w5_rdata[351:344];
  assign w5_45_rdata = w5_rdata[359:352];
  assign w5_46_rdata = w5_rdata[367:360];
  assign w5_47_rdata = w5_rdata[375:368];
  assign w5_48_rdata = w5_rdata[383:376];
  assign w5_49_rdata = w5_rdata[391:384];
  assign w5_50_rdata = w5_rdata[399:392];
  assign w5_51_rdata = w5_rdata[407:400];
  assign w5_52_rdata = w5_rdata[415:408];
  assign w5_53_rdata = w5_rdata[423:416];
  assign w5_54_rdata = w5_rdata[431:424];
  assign w5_55_rdata = w5_rdata[439:432];
  assign w5_56_rdata = w5_rdata[447:440];
  assign w5_57_rdata = w5_rdata[455:448];
  assign w5_58_rdata = w5_rdata[463:456];
  assign w5_59_rdata = w5_rdata[471:464];
  assign w5_60_rdata = w5_rdata[479:472];
  assign w5_61_rdata = w5_rdata[487:480];
  assign w5_62_rdata = w5_rdata[495:488];
  assign w5_63_rdata = w5_rdata[503:496];
  assign w5_64_rdata = w5_rdata[511:504];
  assign w5_65_rdata = w5_rdata[519:512];
  assign w5_66_rdata = w5_rdata[527:520];
  assign w5_67_rdata = w5_rdata[535:528];
  assign w5_68_rdata = w5_rdata[543:536];
  assign w5_69_rdata = w5_rdata[551:544];
  assign w5_70_rdata = w5_rdata[559:552];
  assign w5_71_rdata = w5_rdata[567:560];
  assign w5_72_rdata = w5_rdata[575:568];
  assign w5_73_rdata = w5_rdata[583:576];
  assign w5_74_rdata = w5_rdata[591:584];
  assign w5_75_rdata = w5_rdata[599:592];
  assign w5_76_rdata = w5_rdata[607:600];
  assign w5_77_rdata = w5_rdata[615:608];
  assign w5_78_rdata = w5_rdata[623:616];
  assign w5_79_rdata = w5_rdata[631:624];
  assign w5_80_rdata = w5_rdata[639:632];
  assign w5_81_rdata = w5_rdata[647:640];
  assign w5_82_rdata = w5_rdata[655:648];
  assign w5_83_rdata = w5_rdata[663:656];
  assign w5_84_rdata = w5_rdata[671:664];
  assign w5_85_rdata = w5_rdata[679:672];
  assign w5_86_rdata = w5_rdata[687:680];
  assign w5_87_rdata = w5_rdata[695:688];
  assign w5_88_rdata = w5_rdata[703:696];
  assign w5_89_rdata = w5_rdata[711:704];
  assign w5_90_rdata = w5_rdata[719:712];
  assign w5_91_rdata = w5_rdata[727:720];
  assign w5_92_rdata = w5_rdata[735:728];
  assign w5_93_rdata = w5_rdata[743:736];
  assign w5_94_rdata = w5_rdata[751:744];
  assign w5_95_rdata = w5_rdata[759:752];
  assign w5_96_rdata = w5_rdata[767:760];
  assign w5_97_rdata = w5_rdata[775:768];
  assign w5_98_rdata = w5_rdata[783:776];
  assign w5_99_rdata = w5_rdata[791:784];
  assign w5_100_rdata = w5_rdata[799:792];
  assign w5_101_rdata = w5_rdata[807:800];
  assign w5_102_rdata = w5_rdata[815:808];
  assign w5_103_rdata = w5_rdata[823:816];
  assign w5_104_rdata = w5_rdata[831:824];
  assign w5_105_rdata = w5_rdata[839:832];
  assign w5_106_rdata = w5_rdata[847:840];
  assign w5_107_rdata = w5_rdata[855:848];
  assign w5_108_rdata = w5_rdata[863:856];
  assign w5_109_rdata = w5_rdata[871:864];
  assign w5_110_rdata = w5_rdata[879:872];
  assign w5_111_rdata = w5_rdata[887:880];
  assign w5_112_rdata = w5_rdata[895:888];
  assign w5_113_rdata = w5_rdata[903:896];
  assign w5_114_rdata = w5_rdata[911:904];
  assign w5_115_rdata = w5_rdata[919:912];
  assign w5_116_rdata = w5_rdata[927:920];
  assign w5_117_rdata = w5_rdata[935:928];
  assign w5_118_rdata = w5_rdata[943:936];
  assign w5_119_rdata = w5_rdata[951:944];
  assign w5_120_rdata = w5_rdata[959:952];



endmodule