//==================================================================================================
//  Filename      : w5_rom.v
//  Created On    : 2018-01-07 22:27:49
//  Last Modified : 2018-01-08 12:08:42
//  Revision      : 
//  Author        : YzTong
//  Company       : UESTC
//  Email         : yztong1994@gmail.com
//
//  Description   : 
//
//
//==================================================================================================
module w5_rom(/*autoport*/
//output
      w5_1_rdata,
      w5_2_rdata,
      w5_3_rdata,
      w5_4_rdata,
      w5_5_rdata,
      w5_6_rdata,
      w5_7_rdata,
      w5_8_rdata,
      w5_9_rdata,
      w5_10_rdata,
      w5_11_rdata,
      w5_12_rdata,
      w5_13_rdata,
      w5_14_rdata,
      w5_15_rdata,
      w5_16_rdata,
      w5_17_rdata,
      w5_18_rdata,
      w5_19_rdata,
      w5_20_rdata,
      w5_21_rdata,
      w5_22_rdata,
      w5_23_rdata,
      w5_24_rdata,
      w5_25_rdata,
      w5_26_rdata,
      w5_27_rdata,
      w5_28_rdata,
      w5_29_rdata,
      w5_30_rdata,
      w5_31_rdata,
      w5_32_rdata,
      w5_33_rdata,
      w5_34_rdata,
      w5_35_rdata,
      w5_36_rdata,
      w5_37_rdata,
      w5_38_rdata,
      w5_39_rdata,
      w5_40_rdata,
      w5_41_rdata,
      w5_42_rdata,
      w5_43_rdata,
      w5_44_rdata,
      w5_45_rdata,
      w5_46_rdata,
      w5_47_rdata,
      w5_48_rdata,
      w5_49_rdata,
      w5_50_rdata,
      w5_51_rdata,
      w5_52_rdata,
      w5_53_rdata,
      w5_54_rdata,
      w5_55_rdata,
      w5_56_rdata,
      w5_57_rdata,
      w5_58_rdata,
      w5_59_rdata,
      w5_60_rdata,
      w5_61_rdata,
      w5_62_rdata,
      w5_63_rdata,
      w5_64_rdata,
      w5_65_rdata,
      w5_66_rdata,
      w5_67_rdata,
      w5_68_rdata,
      w5_69_rdata,
      w5_70_rdata,
      w5_71_rdata,
      w5_72_rdata,
      w5_73_rdata,
      w5_74_rdata,
      w5_75_rdata,
      w5_76_rdata,
      w5_77_rdata,
      w5_78_rdata,
      w5_79_rdata,
      w5_80_rdata,
      w5_81_rdata,
      w5_82_rdata,
      w5_83_rdata,
      w5_84_rdata,
      w5_85_rdata,
      w5_86_rdata,
      w5_87_rdata,
      w5_88_rdata,
      w5_89_rdata,
      w5_90_rdata,
      w5_91_rdata,
      w5_92_rdata,
      w5_93_rdata,
      w5_94_rdata,
      w5_95_rdata,
      w5_96_rdata,
      w5_97_rdata,
      w5_98_rdata,
      w5_99_rdata,
      w5_100_rdata,
      w5_101_rdata,
      w5_102_rdata,
      w5_103_rdata,
      w5_104_rdata,
      w5_105_rdata,
      w5_106_rdata,
      w5_107_rdata,
      w5_108_rdata,
      w5_109_rdata,
      w5_110_rdata,
      w5_111_rdata,
      w5_112_rdata,
      w5_113_rdata,
      w5_114_rdata,
      w5_115_rdata,
      w5_116_rdata,
      w5_117_rdata,
      w5_118_rdata,
      w5_119_rdata,
      w5_120_rdata,
//input
      clk,
      w5_raddr);
	
	input clk;
	input [8:0] w5_raddr;
	output[7:0] w5_1_rdata;	
	output[7:0] w5_2_rdata;
	output[7:0] w5_3_rdata;
	output[7:0] w5_4_rdata;
	output[7:0] w5_5_rdata;
	output[7:0] w5_6_rdata;
	output[7:0] w5_7_rdata;
	output[7:0] w5_8_rdata;
	output[7:0] w5_9_rdata;
	output[7:0] w5_10_rdata;
	output[7:0] w5_11_rdata;
	output[7:0] w5_12_rdata;
	output[7:0] w5_13_rdata;
	output[7:0] w5_14_rdata;
	output[7:0] w5_15_rdata;
	output[7:0] w5_16_rdata;
	output[7:0] w5_17_rdata;
	output[7:0] w5_18_rdata;
	output[7:0] w5_19_rdata;
	output[7:0] w5_20_rdata;
	output[7:0] w5_21_rdata;
	output[7:0] w5_22_rdata;
	output[7:0] w5_23_rdata;
	output[7:0] w5_24_rdata;
	output[7:0] w5_25_rdata;
	output[7:0] w5_26_rdata;
	output[7:0] w5_27_rdata;
	output[7:0] w5_28_rdata;
	output[7:0] w5_29_rdata;
	output[7:0] w5_30_rdata;
	output[7:0] w5_31_rdata;
	output[7:0] w5_32_rdata;
	output[7:0] w5_33_rdata;
	output[7:0] w5_34_rdata;
	output[7:0] w5_35_rdata;
	output[7:0] w5_36_rdata;
	output[7:0] w5_37_rdata;
	output[7:0] w5_38_rdata;
	output[7:0] w5_39_rdata;
	output[7:0] w5_40_rdata;
	output[7:0] w5_41_rdata;
	output[7:0] w5_42_rdata;
	output[7:0] w5_43_rdata;
	output[7:0] w5_44_rdata;
	output[7:0] w5_45_rdata;
	output[7:0] w5_46_rdata;
	output[7:0] w5_47_rdata;
	output[7:0] w5_48_rdata;
	output[7:0] w5_49_rdata;
	output[7:0] w5_50_rdata;
	output[7:0] w5_51_rdata;
	output[7:0] w5_52_rdata;
	output[7:0] w5_53_rdata;
	output[7:0] w5_54_rdata;
	output[7:0] w5_55_rdata;
	output[7:0] w5_56_rdata;
	output[7:0] w5_57_rdata;
	output[7:0] w5_58_rdata;
	output[7:0] w5_59_rdata;
	output[7:0] w5_60_rdata;
	output[7:0] w5_61_rdata;
	output[7:0] w5_62_rdata;
	output[7:0] w5_63_rdata;
	output[7:0] w5_64_rdata;
	output[7:0] w5_65_rdata;
	output[7:0] w5_66_rdata;
	output[7:0] w5_67_rdata;
	output[7:0] w5_68_rdata;
	output[7:0] w5_69_rdata;
	output[7:0] w5_70_rdata;
	output[7:0] w5_71_rdata;
	output[7:0] w5_72_rdata;
	output[7:0] w5_73_rdata;
	output[7:0] w5_74_rdata;
	output[7:0] w5_75_rdata;
	output[7:0] w5_76_rdata;
	output[7:0] w5_77_rdata;
	output[7:0] w5_78_rdata;
	output[7:0] w5_79_rdata;
	output[7:0] w5_80_rdata;
	output[7:0] w5_81_rdata;
	output[7:0] w5_82_rdata;
	output[7:0] w5_83_rdata;
	output[7:0] w5_84_rdata;
	output[7:0] w5_85_rdata;
	output[7:0] w5_86_rdata;
	output[7:0] w5_87_rdata;
	output[7:0] w5_88_rdata;
	output[7:0] w5_89_rdata;
	output[7:0] w5_90_rdata;
	output[7:0] w5_91_rdata;
	output[7:0] w5_92_rdata;
	output[7:0] w5_93_rdata;
	output[7:0] w5_94_rdata;
	output[7:0] w5_95_rdata;
	output[7:0] w5_96_rdata;
	output[7:0] w5_97_rdata;
	output[7:0] w5_98_rdata;
	output[7:0] w5_99_rdata;
	output[7:0] w5_100_rdata;
	output[7:0] w5_101_rdata;
	output[7:0] w5_102_rdata;
	output[7:0] w5_103_rdata;
	output[7:0] w5_104_rdata;
	output[7:0] w5_105_rdata;
	output[7:0] w5_106_rdata;
	output[7:0] w5_107_rdata;
	output[7:0] w5_108_rdata;
	output[7:0] w5_109_rdata;
	output[7:0] w5_110_rdata;
	output[7:0] w5_111_rdata;
	output[7:0] w5_112_rdata;
	output[7:0] w5_113_rdata;
	output[7:0] w5_114_rdata;
	output[7:0] w5_115_rdata;
	output[7:0] w5_116_rdata;
	output[7:0] w5_117_rdata;
	output[7:0] w5_118_rdata;
	output[7:0] w5_119_rdata;
	output[7:0] w5_120_rdata;

blk_mem_gen_w5_1_rom w5_1 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_1_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_2_rom w5_2 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_2_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_3_rom w5_3 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_3_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_4_rom w5_4 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_4_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_5_rom w5_5 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_5_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_6_rom w5_6 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_6_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_7_rom w5_7 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_7_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_8_rom w5_8 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_8_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_9_rom w5_9 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_9_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_10_rom w5_10 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_10_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_11_rom w5_11 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_11_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_12_rom w5_12 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_12_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_13_rom w5_13 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_13_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_14_rom w5_14 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_14_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_15_rom w5_15 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_15_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_16_rom w5_16 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_16_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_17_rom w5_17 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_17_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_18_rom w5_18 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_18_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_19_rom w5_19 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_19_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_20_rom w5_20 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_20_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_21_rom w5_21 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_21_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_22_rom w5_22 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_22_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_23_rom w5_23 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_23_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_24_rom w5_24 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_24_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_25_rom w5_25 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_25_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_26_rom w5_26 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_26_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_27_rom w5_27 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_27_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_28_rom w5_28 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_28_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_29_rom w5_29 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_29_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_30_rom w5_30 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_30_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_31_rom w5_31 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_31_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_32_rom w5_32 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_32_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_33_rom w5_33 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_33_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_34_rom w5_34 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_34_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_35_rom w5_35 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_35_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_36_rom w5_36 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_36_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_37_rom w5_37 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_37_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_38_rom w5_38 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_38_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_39_rom w5_39 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_39_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_40_rom w5_40 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_40_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_41_rom w5_41 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_41_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_42_rom w5_42 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_42_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_43_rom w5_43 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_43_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_44_rom w5_44 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_44_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_45_rom w5_45 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_45_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_46_rom w5_46 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_46_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_47_rom w5_47 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_47_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_48_rom w5_48 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_48_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_49_rom w5_49 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_49_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_50_rom w5_50 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_50_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_51_rom w5_51 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_51_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_52_rom w5_52 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_52_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_53_rom w5_53 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_53_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_54_rom w5_54 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_54_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_55_rom w5_55 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_55_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_56_rom w5_56 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_56_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_57_rom w5_57 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_57_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_58_rom w5_58 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_58_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_59_rom w5_59 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_59_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_60_rom w5_60 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_60_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_61_rom w5_61 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_61_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_62_rom w5_62 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_62_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_63_rom w5_63 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_63_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_64_rom w5_64 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_64_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_65_rom w5_65 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_65_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_66_rom w5_66 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_66_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_67_rom w5_67 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_67_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_68_rom w5_68 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_68_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_69_rom w5_69 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_69_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_70_rom w5_70 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_70_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_71_rom w5_71 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_71_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_72_rom w5_72 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_72_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_73_rom w5_73 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_73_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_74_rom w5_74 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_74_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_75_rom w5_75 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_75_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_76_rom w5_76 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_76_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_77_rom w5_77 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_77_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_78_rom w5_78 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_78_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_79_rom w5_79 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_79_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_80_rom w5_80 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_80_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_81_rom w5_81 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_81_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_82_rom w5_82 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_82_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_83_rom w5_83 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_83_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_84_rom w5_84 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_84_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_85_rom w5_85 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_85_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_86_rom w5_86 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_86_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_87_rom w5_87 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_87_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_88_rom w5_88 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_88_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_89_rom w5_89 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_89_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_90_rom w5_90 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_90_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_91_rom w5_91 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_91_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_92_rom w5_92 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_92_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_93_rom w5_93 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_93_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_94_rom w5_94 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_94_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_95_rom w5_95 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_95_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_96_rom w5_96 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_96_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_97_rom w5_97 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_97_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_98_rom w5_98 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_98_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_99_rom w5_99 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_99_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_100_rom w5_100 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_100_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_101_rom w5_101 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_101_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_102_rom w5_102 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_102_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_103_rom w5_103 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_103_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_104_rom w5_104 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_104_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_105_rom w5_105 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_105_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_106_rom w5_106 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_106_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_107_rom w5_107 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_107_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_108_rom w5_108 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_108_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_109_rom w5_109 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_109_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_110_rom w5_110 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_110_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_111_rom w5_111 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_111_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_112_rom w5_112 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_112_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_113_rom w5_113 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_113_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_114_rom w5_114 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_114_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_115_rom w5_115 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_115_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_116_rom w5_116 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_116_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_117_rom w5_117 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_117_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_118_rom w5_118 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_118_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_119_rom w5_119 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_119_rdata)  // output wire [7 : 0] douta
);
blk_mem_gen_w5_120_rom w5_120 (
  .clka(clk),    // input wire clka
  .addra(w5_raddr),  // input wire [8 : 0] addra
  .douta(w5_120_rdata)  // output wire [7 : 0] douta
);




endmodule